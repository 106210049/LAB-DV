package fifo_pkg;
 `include "transaction.sv"
 `include "generator.sv"
 `include "driver.sv"
 `include "monitor.sv"
 `include "scoreboard.sv"
 `include "agent.sv"
 `include "env.sv"
endpackage: fifo_pkg

